`ifndef __USER_EXTERNS_SVH__
`define __USER_EXTERNS_SVH__

`define ENABLED_USER_EXTERNS

`endif // __USER_EXTERNS_SVH__
